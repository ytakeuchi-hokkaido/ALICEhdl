library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity D_ffs is	

  generic(
    In_width : natural := 10;
    sel_width : natural := 2;
    SUM_width : natural := 18;
    cont_width: natural := 9;
    contri_width:natural := 9;
    average_width:natural := 12;
    LT_add_width : natural := 4;
    Add_width: natural := 13
    );

  

  port(
    Clock											:in std_logic;
    In_1, In_2, In_3, In_4, In_5, In_6, In_7, In_8, In_9, In_10 				:in  unsigned((In_width-1) downto 0);
    In_11, In_12, In_13, In_14, In_15, In_16, In_17, In_18, In_19, In_20 			:in  unsigned((In_width-1) downto 0);
    In_21, In_22, In_23, In_24, In_25, In_26, In_27, In_28, In_29, In_30 			:in  unsigned((In_width-1) downto 0);
    In_31, In_32, In_33, In_34, In_35, In_36, In_37, In_38, In_39, In_40 			:in  unsigned((In_width-1) downto 0);
    In_41, In_42, In_43, In_44, In_45, In_46, In_47, In_48, In_49, In_50			:in  unsigned((In_width-1) downto 0); 
    In_51, In_52, In_53, In_54, In_55, In_56, In_57, In_58, In_59, In_60 			:in  unsigned((In_width-1) downto 0);
    In_61, In_62, In_63, In_64, In_65, In_66, In_67, In_68, In_69, In_70 			:in  unsigned((In_width-1) downto 0);
    In_71, In_72, In_73, In_74, In_75, In_76, In_77, In_78, In_79, In_80 			:in  unsigned((In_width-1) downto 0);
    In_81, In_82, In_83, In_84, In_85, In_86, In_87, In_88, In_89, In_90 			:in  unsigned((In_width-1) downto 0);
    In_91, In_92, In_93, In_94, In_95, In_96, In_97, In_98, In_99, In_100 			:in  unsigned((In_width-1) downto 0);
    In_101, In_102, In_103, In_104, In_105, In_106, In_107, In_108, In_109, In_110	        :in  unsigned((In_width-1) downto 0); 
    In_111, In_112, In_113, In_114, In_115, In_116, In_117, In_118, In_119, In_120 	        :in  unsigned((In_width-1) downto 0);
    In_121, In_122, In_123, In_124, In_125, In_126, In_127, In_128, In_129, In_130 	        :in  unsigned((In_width-1) downto 0);
    In_131, In_132, In_133, In_134, In_135, In_136, In_137, In_138, In_139, In_140 	        :in  unsigned((In_width-1) downto 0);
    In_141, In_142, In_143, In_144, In_145, In_146, In_147, In_148, In_149, In_150 	        :in  unsigned((In_width-1) downto 0);
    In_151, In_152, In_153, In_154, In_155, In_156, In_157, In_158, In_159, In_160 	        :in  unsigned((In_width-1) downto 0);
    In_161, In_162, In_163, In_164, In_165, In_166, In_167, In_168, In_169, In_170 	        :in  unsigned((In_width-1) downto 0);
    In_171, In_172, In_173, In_174, In_175, In_176, In_177, In_178, In_179, In_180 	        :in  unsigned((In_width-1) downto 0);
    In_181, In_182, In_183, In_184, In_185, In_186, In_187, In_188, In_189, In_190 	        :in  unsigned((In_width-1) downto 0);
    In_191, In_192, In_193, In_194, In_195, In_196, In_197, In_198, In_199, In_200 	        :in  unsigned((In_width-1) downto 0);
    Df_o1, Df_o2, Df_o3, Df_o4, Df_o5, Df_o6, Df_o7, Df_o8, Df_o9, Df_o10 			:out  unsigned((In_width-1) downto 0);
    Df_o11, Df_o12, Df_o13, Df_o14, Df_o15, Df_o16, Df_o17, Df_o18, Df_o19, Df_o20 		:out  unsigned((In_width-1) downto 0);
    Df_o21, Df_o22, Df_o23, Df_o24, Df_o25, Df_o26, Df_o27, Df_o28, Df_o29, Df_o30 		:out  unsigned((In_width-1) downto 0);
    Df_o31, Df_o32, Df_o33, Df_o34, Df_o35, Df_o36, Df_o37, Df_o38, Df_o39, Df_o40 		:out  unsigned((In_width-1) downto 0);
    Df_o41, Df_o42, Df_o43, Df_o44, Df_o45, Df_o46, Df_o47, Df_o48, Df_o49, Df_o50		:out  unsigned((In_width-1) downto 0); 
    Df_o51, Df_o52, Df_o53, Df_o54, Df_o55, Df_o56, Df_o57, Df_o58, Df_o59, Df_o60 		:out  unsigned((In_width-1) downto 0);
    Df_o61, Df_o62, Df_o63, Df_o64, Df_o65, Df_o66, Df_o67, Df_o68, Df_o69, Df_o70 		:out  unsigned((In_width-1) downto 0);
    Df_o71, Df_o72, Df_o73, Df_o74, Df_o75, Df_o76, Df_o77, Df_o78, Df_o79, Df_o80 		:out  unsigned((In_width-1) downto 0);
    Df_o81, Df_o82, Df_o83, Df_o84, Df_o85, Df_o86, Df_o87, Df_o88, Df_o89, Df_o90 		:out  unsigned((In_width-1) downto 0);
    Df_o91, Df_o92, Df_o93, Df_o94, Df_o95, Df_o96, Df_o97, Df_o98, Df_o99, Df_o100 	:out  unsigned((In_width-1) downto 0);
    Df_o101, Df_o102, Df_o103, Df_o104, Df_o105, Df_o106, Df_o107, Df_o108, Df_o109, Df_o110:out  unsigned((In_width-1) downto 0); 
    Df_o111, Df_o112, Df_o113, Df_o114, Df_o115, Df_o116, Df_o117, Df_o118, Df_o119, Df_o120:out  unsigned((In_width-1) downto 0);
    Df_o121, Df_o122, Df_o123, Df_o124, Df_o125, Df_o126, Df_o127, Df_o128, Df_o129, Df_o130:out  unsigned((In_width-1) downto 0);
    Df_o131, Df_o132, Df_o133, Df_o134, Df_o135, Df_o136, Df_o137, Df_o138, Df_o139, Df_o140:out  unsigned((In_width-1) downto 0);
    Df_o141, Df_o142, Df_o143, Df_o144, Df_o145, Df_o146, Df_o147, Df_o148, Df_o149, Df_o150:out  unsigned((In_width-1) downto 0);
    Df_o151, Df_o152, Df_o153, Df_o154, Df_o155, Df_o156, Df_o157, Df_o158, Df_o159, Df_o160:out  unsigned((In_width-1) downto 0);
    Df_o161, Df_o162, Df_o163, Df_o164, Df_o165, Df_o166, Df_o167, Df_o168, Df_o169, Df_o170:out  unsigned((In_width-1) downto 0);
    Df_o171, Df_o172, Df_o173, Df_o174, Df_o175, Df_o176, Df_o177, Df_o178, Df_o179, Df_o180:out  unsigned((In_width-1) downto 0);
    Df_o181, Df_o182, Df_o183, Df_o184, Df_o185, Df_o186, Df_o187, Df_o188, Df_o189, Df_o190:out  unsigned((In_width-1) downto 0);
    Df_o191, Df_o192, Df_o193, Df_o194, Df_o195, Df_o196, Df_o197, Df_o198, Df_o199, Df_o200:out  unsigned((In_width-1) downto 0)
    );
  
end entity;

architecture rtl of D_ffs is
-- D-flip flop

  component D_ff port(
    Clock :in std_logic;
    Input :in unsigned((In_width-1) downto 0):= "0000000000";
    Output :out unsigned((In_width-1) downto 0):= "0000000000"
    );
end component;
-- D-flip flop
begin
  D_ff1:D_ff port map(Clock => Clock, Input => In_1, Output => Df_o1);
  D_ff2:D_ff port map(Clock => Clock, Input => In_2, Output => Df_o2);
  D_ff3:D_ff port map(Clock => Clock, Input => In_3, Output => Df_o3);
  D_ff4:D_ff port map(Clock => Clock, Input => In_4, Output => Df_o4);
  D_ff5:D_ff port map(Clock => Clock, Input => In_5, Output => Df_o5);
  D_ff6:D_ff port map(Clock => Clock, Input => In_6, Output => Df_o6);
  D_ff7:D_ff port map(Clock => Clock, Input => In_7, Output => Df_o7);
  D_ff8:D_ff port map(Clock => Clock, Input => In_8, Output => Df_o8);
  D_ff9:D_ff port map(Clock => Clock, Input => In_9, Output => Df_o9);
  D_ff10:D_ff port map(Clock => Clock, Input => In_10, Output => Df_o10);
  D_ff11:D_ff port map(Clock => Clock, Input => In_11, Output => Df_o11);
  D_ff12:D_ff port map(Clock => Clock, Input => In_12, Output => Df_o12);
  D_ff13:D_ff port map(Clock => Clock, Input => In_13, Output => Df_o13);
  D_ff14:D_ff port map(Clock => Clock, Input => In_14, Output => Df_o14);
  D_ff15:D_ff port map(Clock => Clock, Input => In_15, Output => Df_o15);
  D_ff16:D_ff port map(Clock => Clock, Input => In_16, Output => Df_o16);
  D_ff17:D_ff port map(Clock => Clock, Input => In_17, Output => Df_o17);
  D_ff18:D_ff port map(Clock => Clock, Input => In_18, Output => Df_o18);
  D_ff19:D_ff port map(Clock => Clock, Input => In_19, Output => Df_o19);
  D_ff20:D_ff port map(Clock => Clock, Input => In_20, Output => Df_o20);
  D_ff21:D_ff port map(Clock => Clock, Input => In_21, Output => Df_o21);
  D_ff22:D_ff port map(Clock => Clock, Input => In_22, Output => Df_o22);
  D_ff23:D_ff port map(Clock => Clock, Input => In_23, Output => Df_o23);
  D_ff24:D_ff port map(Clock => Clock, Input => In_24, Output => Df_o24);
  D_ff25:D_ff port map(Clock => Clock, Input => In_25, Output => Df_o25);
  D_ff26:D_ff port map(Clock => Clock, Input => In_26, Output => Df_o26);
  D_ff27:D_ff port map(Clock => Clock, Input => In_27, Output => Df_o27);
  D_ff28:D_ff port map(Clock => Clock, Input => In_28, Output => Df_o28);
  D_ff29:D_ff port map(Clock => Clock, Input => In_29, Output => Df_o29);
  D_ff30:D_ff port map(Clock => Clock, Input => In_30, Output => Df_o30);
  D_ff31:D_ff port map(Clock => Clock, Input => In_31, Output => Df_o31);
  D_ff32:D_ff port map(Clock => Clock, Input => In_32, Output => Df_o32);
  D_ff33:D_ff port map(Clock => Clock, Input => In_33, Output => Df_o33);
  D_ff34:D_ff port map(Clock => Clock, Input => In_34, Output => Df_o34);
  D_ff35:D_ff port map(Clock => Clock, Input => In_35, Output => Df_o35);
  D_ff36:D_ff port map(Clock => Clock, Input => In_36, Output => Df_o36);
  D_ff37:D_ff port map(Clock => Clock, Input => In_37, Output => Df_o37);
  D_ff38:D_ff port map(Clock => Clock, Input => In_38, Output => Df_o38);
  D_ff39:D_ff port map(Clock => Clock, Input => In_39, Output => Df_o39);
  D_ff40:D_ff port map(Clock => Clock, Input => In_40, Output => Df_o40);
  D_ff41:D_ff port map(Clock => Clock, Input => In_41, Output => Df_o41);
  D_ff42:D_ff port map(Clock => Clock, Input => In_42, Output => Df_o42);
  D_ff43:D_ff port map(Clock => Clock, Input => In_43, Output => Df_o43);
  D_ff44:D_ff port map(Clock => Clock, Input => In_44, Output => Df_o44);
  D_ff45:D_ff port map(Clock => Clock, Input => In_45, Output => Df_o45);
  D_ff46:D_ff port map(Clock => Clock, Input => In_46, Output => Df_o46);
  D_ff47:D_ff port map(Clock => Clock, Input => In_47, Output => Df_o47);
  D_ff48:D_ff port map(Clock => Clock, Input => In_48, Output => Df_o48);
  D_ff49:D_ff port map(Clock => Clock, Input => In_49, Output => Df_o49);
  D_ff50:D_ff port map(Clock => Clock, Input => In_50, Output => Df_o50);
  D_ff51:D_ff port map(Clock => Clock, Input => In_51, Output => Df_o51);
  D_ff52:D_ff port map(Clock => Clock, Input => In_52, Output => Df_o52);
  D_ff53:D_ff port map(Clock => Clock, Input => In_53, Output => Df_o53);
  D_ff54:D_ff port map(Clock => Clock, Input => In_54, Output => Df_o54);
  D_ff55:D_ff port map(Clock => Clock, Input => In_55, Output => Df_o55);
  D_ff56:D_ff port map(Clock => Clock, Input => In_56, Output => Df_o56);
  D_ff57:D_ff port map(Clock => Clock, Input => In_57, Output => Df_o57);
  D_ff58:D_ff port map(Clock => Clock, Input => In_58, Output => Df_o58);
  D_ff59:D_ff port map(Clock => Clock, Input => In_59, Output => Df_o59);
  D_ff60:D_ff port map(Clock => Clock, Input => In_60, Output => Df_o60);
  D_ff61:D_ff port map(Clock => Clock, Input => In_61, Output => Df_o61);
  D_ff62:D_ff port map(Clock => Clock, Input => In_62, Output => Df_o62);
  D_ff63:D_ff port map(Clock => Clock, Input => In_63, Output => Df_o63);
  D_ff64:D_ff port map(Clock => Clock, Input => In_64, Output => Df_o64);
  D_ff65:D_ff port map(Clock => Clock, Input => In_65, Output => Df_o65);
  D_ff66:D_ff port map(Clock => Clock, Input => In_66, Output => Df_o66);
  D_ff67:D_ff port map(Clock => Clock, Input => In_67, Output => Df_o67);
  D_ff68:D_ff port map(Clock => Clock, Input => In_68, Output => Df_o68);
  D_ff69:D_ff port map(Clock => Clock, Input => In_69, Output => Df_o69);
  D_ff70:D_ff port map(Clock => Clock, Input => In_70, Output => Df_o70);
  D_ff71:D_ff port map(Clock => Clock, Input => In_71, Output => Df_o71);
  D_ff72:D_ff port map(Clock => Clock, Input => In_72, Output => Df_o72);
  D_ff73:D_ff port map(Clock => Clock, Input => In_73, Output => Df_o73);
  D_ff74:D_ff port map(Clock => Clock, Input => In_74, Output => Df_o74);
  D_ff75:D_ff port map(Clock => Clock, Input => In_75, Output => Df_o75);
  D_ff76:D_ff port map(Clock => Clock, Input => In_76, Output => Df_o76);
  D_ff77:D_ff port map(Clock => Clock, Input => In_77, Output => Df_o77);
  D_ff78:D_ff port map(Clock => Clock, Input => In_78, Output => Df_o78);
  D_ff79:D_ff port map(Clock => Clock, Input => In_79, Output => Df_o79);
  D_ff80:D_ff port map(Clock => Clock, Input => In_80, Output => Df_o80);
  D_ff81:D_ff port map(Clock => Clock, Input => In_81, Output => Df_o81);
  D_ff82:D_ff port map(Clock => Clock, Input => In_82, Output => Df_o82);
  D_ff83:D_ff port map(Clock => Clock, Input => In_83, Output => Df_o83);
  D_ff84:D_ff port map(Clock => Clock, Input => In_84, Output => Df_o84);
  D_ff85:D_ff port map(Clock => Clock, Input => In_85, Output => Df_o85);
  D_ff86:D_ff port map(Clock => Clock, Input => In_86, Output => Df_o86);
  D_ff87:D_ff port map(Clock => Clock, Input => In_87, Output => Df_o87);
  D_ff88:D_ff port map(Clock => Clock, Input => In_88, Output => Df_o88);
  D_ff89:D_ff port map(Clock => Clock, Input => In_89, Output => Df_o89);
  D_ff90:D_ff port map(Clock => Clock, Input => In_90, Output => Df_o90);
  D_ff91:D_ff port map(Clock => Clock, Input => In_91, Output => Df_o91);
  D_ff92:D_ff port map(Clock => Clock, Input => In_92, Output => Df_o92);
  D_ff93:D_ff port map(Clock => Clock, Input => In_93, Output => Df_o93);
  D_ff94:D_ff port map(Clock => Clock, Input => In_94, Output => Df_o94);
  D_ff95:D_ff port map(Clock => Clock, Input => In_95, Output => Df_o95);
  D_ff96:D_ff port map(Clock => Clock, Input => In_96, Output => Df_o96);
  D_ff97:D_ff port map(Clock => Clock, Input => In_97, Output => Df_o97);
  D_ff98:D_ff port map(Clock => Clock, Input => In_98, Output => Df_o98);
  D_ff99:D_ff port map(Clock => Clock, Input => In_99, Output => Df_o99);
  D_ff100:D_ff port map(Clock => Clock, Input => In_100, Output => Df_o100);
  D_ff101:D_ff port map(Clock => Clock, Input => In_101, Output => Df_o101);
  D_ff102:D_ff port map(Clock => Clock, Input => In_102, Output => Df_o102);
  D_ff103:D_ff port map(Clock => Clock, Input => In_103, Output => Df_o103);
  D_ff104:D_ff port map(Clock => Clock, Input => In_104, Output => Df_o104);
  D_ff105:D_ff port map(Clock => Clock, Input => In_105, Output => Df_o105);
  D_ff106:D_ff port map(Clock => Clock, Input => In_106, Output => Df_o106);
  D_ff107:D_ff port map(Clock => Clock, Input => In_107, Output => Df_o107);
  D_ff108:D_ff port map(Clock => Clock, Input => In_108, Output => Df_o108);
  D_ff109:D_ff port map(Clock => Clock, Input => In_109, Output => Df_o109);
  D_ff110:D_ff port map(Clock => Clock, Input => In_110, Output => Df_o110);
  D_ff111:D_ff port map(Clock => Clock, Input => In_111, Output => Df_o111);
  D_ff112:D_ff port map(Clock => Clock, Input => In_112, Output => Df_o112);
  D_ff113:D_ff port map(Clock => Clock, Input => In_113, Output => Df_o113);
  D_ff114:D_ff port map(Clock => Clock, Input => In_114, Output => Df_o114);
  D_ff115:D_ff port map(Clock => Clock, Input => In_115, Output => Df_o115);
  D_ff116:D_ff port map(Clock => Clock, Input => In_116, Output => Df_o116);
  D_ff117:D_ff port map(Clock => Clock, Input => In_117, Output => Df_o117);
  D_ff118:D_ff port map(Clock => Clock, Input => In_118, Output => Df_o118);
  D_ff119:D_ff port map(Clock => Clock, Input => In_119, Output => Df_o119);
  D_ff120:D_ff port map(Clock => Clock, Input => In_120, Output => Df_o120);
  D_ff121:D_ff port map(Clock => Clock, Input => In_121, Output => Df_o121);
  D_ff122:D_ff port map(Clock => Clock, Input => In_122, Output => Df_o122);
  D_ff123:D_ff port map(Clock => Clock, Input => In_123, Output => Df_o123);
  D_ff124:D_ff port map(Clock => Clock, Input => In_124, Output => Df_o124);
  D_ff125:D_ff port map(Clock => Clock, Input => In_125, Output => Df_o125);
  D_ff126:D_ff port map(Clock => Clock, Input => In_126, Output => Df_o126);
  D_ff127:D_ff port map(Clock => Clock, Input => In_127, Output => Df_o127);
  D_ff128:D_ff port map(Clock => Clock, Input => In_128, Output => Df_o128);
  D_ff129:D_ff port map(Clock => Clock, Input => In_129, Output => Df_o129);
  D_ff130:D_ff port map(Clock => Clock, Input => In_130, Output => Df_o130);
  D_ff131:D_ff port map(Clock => Clock, Input => In_131, Output => Df_o131);
  D_ff132:D_ff port map(Clock => Clock, Input => In_132, Output => Df_o132);
  D_ff133:D_ff port map(Clock => Clock, Input => In_133, Output => Df_o133);
  D_ff134:D_ff port map(Clock => Clock, Input => In_134, Output => Df_o134);
  D_ff135:D_ff port map(Clock => Clock, Input => In_135, Output => Df_o135);
  D_ff136:D_ff port map(Clock => Clock, Input => In_136, Output => Df_o136);
  D_ff137:D_ff port map(Clock => Clock, Input => In_137, Output => Df_o137);
  D_ff138:D_ff port map(Clock => Clock, Input => In_138, Output => Df_o138);
  D_ff139:D_ff port map(Clock => Clock, Input => In_139, Output => Df_o139);
  D_ff140:D_ff port map(Clock => Clock, Input => In_140, Output => Df_o140);
  D_ff141:D_ff port map(Clock => Clock, Input => In_141, Output => Df_o141);
  D_ff142:D_ff port map(Clock => Clock, Input => In_142, Output => Df_o142);
  D_ff143:D_ff port map(Clock => Clock, Input => In_143, Output => Df_o143);
  D_ff144:D_ff port map(Clock => Clock, Input => In_144, Output => Df_o144);
  D_ff145:D_ff port map(Clock => Clock, Input => In_145, Output => Df_o145);
  D_ff146:D_ff port map(Clock => Clock, Input => In_146, Output => Df_o146);
  D_ff147:D_ff port map(Clock => Clock, Input => In_147, Output => Df_o147);
  D_ff148:D_ff port map(Clock => Clock, Input => In_148, Output => Df_o148);
  D_ff149:D_ff port map(Clock => Clock, Input => In_149, Output => Df_o149);
  D_ff150:D_ff port map(Clock => Clock, Input => In_150, Output => Df_o150);
  D_ff151:D_ff port map(Clock => Clock, Input => In_151, Output => Df_o151);
  D_ff152:D_ff port map(Clock => Clock, Input => In_152, Output => Df_o152);
  D_ff153:D_ff port map(Clock => Clock, Input => In_153, Output => Df_o153);
  D_ff154:D_ff port map(Clock => Clock, Input => In_154, Output => Df_o154);
  D_ff155:D_ff port map(Clock => Clock, Input => In_155, Output => Df_o155);
  D_ff156:D_ff port map(Clock => Clock, Input => In_156, Output => Df_o156);
  D_ff157:D_ff port map(Clock => Clock, Input => In_157, Output => Df_o157);
  D_ff158:D_ff port map(Clock => Clock, Input => In_158, Output => Df_o158);
  D_ff159:D_ff port map(Clock => Clock, Input => In_159, Output => Df_o159);
  D_ff160:D_ff port map(Clock => Clock, Input => In_160, Output => Df_o160);
  D_ff161:D_ff port map(Clock => Clock, Input => In_161, Output => Df_o161);
  D_ff162:D_ff port map(Clock => Clock, Input => In_162, Output => Df_o162);
  D_ff163:D_ff port map(Clock => Clock, Input => In_163, Output => Df_o163);
  D_ff164:D_ff port map(Clock => Clock, Input => In_164, Output => Df_o164);
  D_ff165:D_ff port map(Clock => Clock, Input => In_165, Output => Df_o165);
  D_ff166:D_ff port map(Clock => Clock, Input => In_166, Output => Df_o166);
  D_ff167:D_ff port map(Clock => Clock, Input => In_167, Output => Df_o167);
  D_ff168:D_ff port map(Clock => Clock, Input => In_168, Output => Df_o168);
  D_ff169:D_ff port map(Clock => Clock, Input => In_169, Output => Df_o169);
  D_ff170:D_ff port map(Clock => Clock, Input => In_170, Output => Df_o170);
  D_ff171:D_ff port map(Clock => Clock, Input => In_171, Output => Df_o171);
  D_ff172:D_ff port map(Clock => Clock, Input => In_172, Output => Df_o172);
  D_ff173:D_ff port map(Clock => Clock, Input => In_173, Output => Df_o173);
  D_ff174:D_ff port map(Clock => Clock, Input => In_174, Output => Df_o174);
  D_ff175:D_ff port map(Clock => Clock, Input => In_175, Output => Df_o175);
  D_ff176:D_ff port map(Clock => Clock, Input => In_176, Output => Df_o176);
  D_ff177:D_ff port map(Clock => Clock, Input => In_177, Output => Df_o177);
  D_ff178:D_ff port map(Clock => Clock, Input => In_178, Output => Df_o178);
  D_ff179:D_ff port map(Clock => Clock, Input => In_179, Output => Df_o179);
  D_ff180:D_ff port map(Clock => Clock, Input => In_180, Output => Df_o180);
  D_ff181:D_ff port map(Clock => Clock, Input => In_181, Output => Df_o181);
  D_ff182:D_ff port map(Clock => Clock, Input => In_182, Output => Df_o182);
  D_ff183:D_ff port map(Clock => Clock, Input => In_183, Output => Df_o183);
  D_ff184:D_ff port map(Clock => Clock, Input => In_184, Output => Df_o184);
  D_ff185:D_ff port map(Clock => Clock, Input => In_185, Output => Df_o185);
  D_ff186:D_ff port map(Clock => Clock, Input => In_186, Output => Df_o186);
  D_ff187:D_ff port map(Clock => Clock, Input => In_187, Output => Df_o187);
  D_ff188:D_ff port map(Clock => Clock, Input => In_188, Output => Df_o188);
  D_ff189:D_ff port map(Clock => Clock, Input => In_189, Output => Df_o189);
  D_ff190:D_ff port map(Clock => Clock, Input => In_190, Output => Df_o190);
  D_ff191:D_ff port map(Clock => Clock, Input => In_191, Output => Df_o191);
  D_ff192:D_ff port map(Clock => Clock, Input => In_192, Output => Df_o192);
  D_ff193:D_ff port map(Clock => Clock, Input => In_193, Output => Df_o193);
  D_ff194:D_ff port map(Clock => Clock, Input => In_194, Output => Df_o194);
  D_ff195:D_ff port map(Clock => Clock, Input => In_195, Output => Df_o195);
  D_ff196:D_ff port map(Clock => Clock, Input => In_196, Output => Df_o196);
  D_ff197:D_ff port map(Clock => Clock, Input => In_197, Output => Df_o197);
  D_ff198:D_ff port map(Clock => Clock, Input => In_198, Output => Df_o198);
  D_ff199:D_ff port map(Clock => Clock, Input => In_199, Output => Df_o199);
  D_ff200:D_ff port map(Clock => Clock, Input => In_200, Output => Df_o200);
end rtl;
